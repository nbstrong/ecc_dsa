library IEEE;
use IEEE.std_logic_1164.all;
--------------------------------------------------------------------------------
entity riscv is
    port (
        clkIn : in    std_logic;
        rstIn : in    std_logic
    );
end riscv;
--------------------------------------------------------------------------------
architecture behav of riscv is
    -- CONSTANTS ---------------------------------------------------------------
    -- SIGNALS -----------------------------------------------------------------
    -- ALIASES -----------------------------------------------------------------
    -- ATTRIBUTES --------------------------------------------------------------
begin
end behav;